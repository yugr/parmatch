module M #(parameter real TCK) ();
endmodule

M #(.TCK(0)) m;

