`ifdef GPIO_ADDRESS
endmodule
`endif /* GPIO_ADDRESS */
