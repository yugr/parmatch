module A #(parameter A, parameter B, parameter C) ();
endmodule

module A #(parameter A, parameter B) ();
endmodule

A #(.A(1)) a;

